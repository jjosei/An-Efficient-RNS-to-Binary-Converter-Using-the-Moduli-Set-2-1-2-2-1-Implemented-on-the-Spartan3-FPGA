library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity sixbitdec is
port(

        input  :in std_logic_vector(8 downto 0);

	    output :out std_logic_vector (20 downto 0)

);
end sixbitdec;


architecture Behavioral of sixbitdec is



begin

    with input select

            output   <= b"000_0001_000_0001_000_0001" when "000000000",

                        b"000_0001_000_0001_100_1111" when "000000001",
                        b"000_0001_000_0001_001_0010" when "000000010",
                        b"000_0001_000_0001_000_0110" when "000000011",
                        b"000_0001_000_0001_100_1100" when "000000100",
                        b"000_0001_000_0001_010_0100" when "000000101",
                        b"000_0001_000_0001_010_0000" when "000000110",
                        b"000_0001_000_0001_000_1111" when "000000111",
                        b"000_0001_000_0001_000_0000" when "000001000",
                        b"000_0001_000_0001_000_0100" when "000001001",

                        b"000_0001_100_1111_000_0001" when "000001010",
                        b"000_0001_100_1111_100_1111" when "000001011",
                        b"000_0001_100_1111_001_0010" when "000001100",
                        b"000_0001_100_1111_000_0110" when "000001101",
                        b"000_0001_100_1111_100_1100" when "000001110",
                        b"000_0001_100_1111_010_0100" when "000001111",
                        b"000_0001_100_1111_010_0000" when "000010000",
                        b"000_0001_100_1111_000_1111" when "000010001",
                        b"000_0001_100_1111_000_0000" when "000010010",
                        b"000_0001_100_1111_000_0100" when "000010011",

                        b"000_0001_001_0010_000_0001" when "000010100",
                        b"000_0001_001_0010_100_1111" when "000010101",
                        b"000_0001_001_0010_001_0010" when "000010110",
                        b"000_0001_001_0010_000_0110" when "000010111",
                        b"000_0001_001_0010_100_1100" when "000011000",
                        b"000_0001_001_0010_010_0100" when "000011001",
                        b"000_0001_001_0010_010_0000" when "000011010",
                        b"000_0001_001_0010_000_1111" when "000011011",
                        b"000_0001_001_0010_000_0000" when "000011100",
                        b"000_0001_001_0010_000_0100" when "000011101",

                        b"000_0001_000_0110_000_0001" when "000011110",
                        b"000_0001_000_0110_100_1111" when "000011111",
                        b"000_0001_000_0110_001_0010" when "000100000",
                        b"000_0001_000_0110_000_0110" when "000100001",
                        b"000_0001_000_0110_100_1100" when "000100010",
                        b"000_0001_000_0110_010_0100" when "000100011",
                        b"000_0001_000_0110_010_0000" when "000100100",
                        b"000_0001_000_0110_000_1111" when "000100101",
                        b"000_0001_000_0110_000_0000" when "000100110",
                        b"000_0001_000_0110_000_0100" when "000100111",

                        b"000_0001_100_1100_000_0001" when "000101000",
                        b"000_0001_100_1100_100_1111" when "000101001",
                        b"000_0001_100_1100_001_0010" when "000101010",
                        b"000_0001_100_1100_000_0110" when "000101011",
                        b"000_0001_100_1100_100_1100" when "000101100",
                        b"000_0001_100_1100_010_0100" when "000101101",
                        b"000_0001_100_1100_010_0000" when "000101110",
                        b"000_0001_100_1100_000_1111" when "000101111",
                        b"000_0001_100_1100_000_0000" when "000110000",
                        b"000_0001_100_1100_000_0100" when "000110001",

                        b"000_0001_010_0100_000_0001" when "000110010",
                        b"000_0001_010_0100_100_1111" when "000110011",
                        b"000_0001_010_0100_001_0010" when "000110100",
                        b"000_0001_010_0100_000_0110" when "000110101",
                        b"000_0001_010_0100_100_1100" when "000110110",
                        b"000_0001_010_0100_010_0100" when "000110111",
                        b"000_0001_010_0100_010_0000" when "000111000",
                        b"000_0001_010_0100_000_1111" when "000111001",
                        b"000_0001_010_0100_000_0000" when "000111010",
                        b"000_0001_010_0100_000_0100" when "000111011",

                        b"000_0001_010_0000_000_0001" when "000111100",
                        b"000_0001_010_0000_100_1111" when "000111101",
                        b"000_0001_010_0000_001_0010" when "000111110",
                        b"000_0001_010_0000_000_0110" when "000111111",
                        b"000_0001_010_0000_100_1100" when "001000000",
                        b"000_0001_010_0000_010_0100" when "001000001",
                        b"000_0001_010_0000_010_0000" when "001000010",
                        b"000_0001_010_0000_000_1111" when "001000011",
                        b"000_0001_010_0000_000_0000" when "001000100",
                        b"000_0001_010_0000_000_0100" when "001000101",

                        b"000_0001_000_1111_000_0001" when "001000110",
                        b"000_0001_000_1111_100_1111" when "001000111",
                        b"000_0001_000_1111_001_0010" when "001001000",
                        b"000_0001_000_1111_000_0110" when "001001001",
                        b"000_0001_000_1111_100_1100" when "001001010",
                        b"000_0001_000_1111_010_0100" when "001001011",
                        b"000_0001_000_1111_010_0000" when "001001100",
                        b"000_0001_000_1111_000_1111" when "001001101",
                        b"000_0001_000_1111_000_0000" when "001001110",
                        b"000_0001_000_1111_000_0100" when "001001111",

                        b"000_0001_000_0000_000_0001" when "001010000",
                        b"000_0001_000_0000_100_1111" when "001010001",
                        b"000_0001_000_0000_001_0010" when "001010010",
                        b"000_0001_000_0000_000_0110" when "001010011",
                        b"000_0001_000_0000_100_1100" when "001010100",
                        b"000_0001_000_0000_010_0100" when "001010101",
                        b"000_0001_000_0000_010_0000" when "001010110",
                        b"000_0001_000_0000_000_1111" when "001010111",
                        b"000_0001_000_0000_000_0000" when "001011000",
                        b"000_0001_000_0000_000_0100" when "001011001",

                        b"000_0001_000_0100_000_0001" when "001011010",
                        b"000_0001_000_0100_100_1111" when "001011011",
                        b"000_0001_000_0100_001_0010" when "001011100",
                        b"000_0001_000_0100_000_0110" when "001011101",
                        b"000_0001_000_0100_100_1100" when "001011110",
                        b"000_0001_000_0100_010_0100" when "001011111",
                        b"000_0001_000_0100_010_0000" when "001100000",
                        b"000_0001_000_0100_000_1111" when "001100001",
                        b"000_0001_000_0100_000_0000" when "001100010",
                        b"000_0001_000_0100_000_0100" when "001100011",

                        b"100_1111_000_0001_000_0001" when "001100100",
                        b"100_1111_000_0001_100_1111" when "001100101",
                        b"100_1111_000_0001_001_0010" when "001100110",
                        b"100_1111_000_0001_000_0110" when "001100111",
                        b"100_1111_000_0001_100_1100" when "001101000",
                        b"100_1111_000_0001_010_0100" when "001101001",
                        b"100_1111_000_0001_010_0000" when "001101010",
                        b"100_1111_000_0001_000_1111" when "001101011",
                        b"100_1111_000_0001_000_0000" when "001101100",
                        b"100_1111_000_0001_000_0100" when "001101101",

                        b"100_1111_100_1111_000_0001" when "001101110",
                        b"100_1111_100_1111_100_1111" when "001101111",
                        b"100_1111_100_1111_001_0010" when "001110000",
                        b"100_1111_100_1111_000_0110" when "001110001",
                        b"100_1111_100_1111_100_1100" when "001110010",
                        b"100_1111_100_1111_010_0100" when "001110011",
                        b"100_1111_100_1111_010_0000" when "001110100",
                        b"100_1111_100_1111_000_1111" when "001110101",
                        b"100_1111_100_1111_000_0000" when "001110110",
                        b"100_1111_100_1111_000_0100" when "001110111",

                        b"100_1111_001_0010_000_0001" when "001111000",
                        b"100_1111_001_0010_100_1111" when "001111001",
                        b"100_1111_001_0010_001_0010" when "001111010",
                        b"100_1111_001_0010_000_0110" when "001111011",
                        b"100_1111_001_0010_100_1100" when "001111100",
                        b"100_1111_001_0010_010_0100" when "001111101",
                        b"100_1111_001_0010_010_0000" when "001111110",
                        b"100_1111_001_0010_000_1111" when "001111111",
                        b"100_1111_001_0010_000_0000" when "010000000",
                        b"100_1111_001_0010_000_0100" when "010000001",

                        b"100_1111_000_0110_000_0001" when "010000010",
                        b"100_1111_000_0110_100_1111" when "010000011",
                        b"100_1111_000_0110_001_0010" when "010000100",
                        b"100_1111_000_0110_000_0110" when "010000101",
                        b"100_1111_000_0110_100_1100" when "010000110",
                        b"100_1111_000_0110_010_0100" when "010000111",
                        b"100_1111_000_0110_010_0000" when "010001000",
                        b"100_1111_000_0110_000_1111" when "010001001",
                        b"100_1111_000_0110_000_0000" when "010001010",
                        b"100_1111_000_0110_000_0100" when "010001011",

                        b"100_1111_100_1100_000_0001" when "010001100",
                        b"100_1111_100_1100_100_1111" when "010001101",
                        b"100_1111_100_1100_001_0010" when "010001110",
                        b"100_1111_100_1100_000_0110" when "010001111",
                        b"100_1111_100_1100_100_1100" when "010010000",
                        b"100_1111_100_1100_010_0100" when "010010001",
                        b"100_1111_100_1100_010_0000" when "010010010",
                        b"100_1111_100_1100_000_1111" when "010010011",
                        b"100_1111_100_1100_000_0000" when "010010100",
                        b"100_1111_100_1100_000_0100" when "010010101",

                        b"100_1111_010_0100_000_0001" when "010010110",
                        b"100_1111_010_0100_100_1111" when "010010111",
                        b"100_1111_010_0100_001_0010" when "010011000",
                        b"100_1111_010_0100_000_0110" when "010011001",
                        b"100_1111_010_0100_100_1100" when "010011010",
                        b"100_1111_010_0100_010_0100" when "010011011",
                        b"100_1111_010_0100_010_0000" when "010011100",
                        b"100_1111_010_0100_000_1111" when "010011101",
                        b"100_1111_010_0100_000_0000" when "010011110",
                        b"100_1111_010_0100_000_0100" when "010011111",
								
                        b"100_1111_010_0000_000_0001" when "010100000",
                        b"100_1111_010_0000_100_1111" when "010100001",
                        b"100_1111_010_0000_001_0010" when "010100010",
                        b"100_1111_010_0000_000_0110" when "010100011",
                        b"100_1111_010_0000_100_1100" when "010100100",
                        b"100_1111_010_0000_010_0100" when "010100101",
                        b"100_1111_010_0000_010_0000" when "010100110",
                        b"100_1111_010_0000_000_1111" when "010100111",
                        b"100_1111_010_0000_000_0000" when "010101000",
                        b"100_1111_010_0000_000_0100" when "010101001",

                        b"100_1111_000_1111_000_0001" when "010101010",
                        b"100_1111_000_1111_100_1111" when "010101011",
                        b"100_1111_000_1111_001_0010" when "010101100",
                        b"100_1111_000_1111_000_0110" when "010101101",
                        b"100_1111_000_1111_100_1100" when "010101110",
                        b"100_1111_000_1111_010_0100" when "010101111",
                        b"100_1111_000_1111_010_0000" when "010110000",
                        b"100_1111_000_1111_000_1111" when "010110001",
                        b"100_1111_000_1111_000_0000" when "010110010",
                        b"100_1111_000_1111_000_0100" when "010110011",

                        b"100_1111_000_0000_000_0001" when "010110100",
                        b"100_1111_000_0000_100_1111" when "010110101",
                        b"100_1111_000_0000_001_0010" when "010110110",
                        b"100_1111_000_0000_000_0110" when "010110111",
                        b"100_1111_000_0000_100_1100" when "010111000",
                        b"100_1111_000_0000_010_0100" when "010111001",
                        b"100_1111_000_0000_010_0000" when "010111010",
                        b"100_1111_000_0000_000_1111" when "010111011",
                        b"100_1111_000_0000_000_0000" when "010111100",
                        b"100_1111_000_0000_000_0100" when "010111101",

                        b"100_1111_000_0100_000_0001" when "010111110",
                        b"100_1111_000_0100_100_1111" when "010111111",
                        b"100_1111_000_0100_001_0010" when "011000000",
                        b"100_1111_000_0100_000_0110" when "011000001",
                        b"100_1111_000_0100_100_1100" when "011000010",
                        b"100_1111_000_0100_010_0100" when "011000011",
                        b"100_1111_000_0100_010_0000" when "011000100",
                        b"100_1111_000_0100_000_1111" when "011000101",
                        b"100_1111_000_0100_000_0000" when "011000110",
                        b"100_1111_000_0100_000_0100" when "011000111",

                        b"001_0010_000_0001_000_0001" when "011001000",
                        b"001_0010_000_0001_100_1111" when "011001001",
                        b"001_0010_000_0001_001_0010" when "011001010",
                        b"001_0010_000_0001_000_0110" when "011001011",
                        b"001_0010_000_0001_100_1100" when "011001100",
                        b"001_0010_000_0001_010_0100" when "011001101",
                        b"001_0010_000_0001_010_0000" when "011001110",
                        b"001_0010_000_0001_000_1111" when "011001111",
                        b"001_0010_000_0001_000_0000" when "011010000",
                        b"001_0010_000_0001_000_0100" when "011010001",

                        b"001_0010_100_1111_000_0001" when "011010010",
                        b"001_0010_100_1111_100_1111" when "011010011",
                        b"001_0010_100_1111_001_0010" when "011010100",
                        b"001_0010_100_1111_000_0110" when "011010101",
                        b"001_0010_100_1111_100_1100" when "011010110",
                        b"001_0010_100_1111_010_0100" when "011010111",
                        b"001_0010_100_1111_010_0000" when "011011000",
                        b"001_0010_100_1111_000_1111" when "011011001",
                        b"001_0010_100_1111_000_0000" when "011011010",
                        b"001_0010_100_1111_000_0100" when "011011011",

                        b"001_0010_001_0010_000_0001" when "011011100",
                        b"001_0010_001_0010_100_1111" when "011011101",
                        b"001_0010_001_0010_001_0010" when "011011110",
                        b"001_0010_001_0010_000_0110" when "011011111",
                        b"001_0010_001_0010_100_1100" when "011100000",
                        b"001_0010_001_0010_010_0100" when "011100001",
                        b"001_0010_001_0010_010_0000" when "011100010",
                        b"001_0010_001_0010_000_1111" when "011100011",
                        b"001_0010_001_0010_000_0000" when "011100100",
                        b"001_0010_001_0010_000_0100" when "011100101",

                        b"001_0010_000_0110_000_0001" when "011100110",
                        b"001_0010_000_0110_100_1111" when "011100111",
                        b"001_0010_000_0110_001_0010" when "011101000",
                        b"001_0010_000_0110_000_0110" when "011101001",
                        b"001_0010_000_0110_100_1100" when "011101010",
                        b"001_0010_000_0110_010_0100" when "011101011",
                        b"001_0010_000_0110_010_0000" when "011101100",
                        b"001_0010_000_0110_000_1111" when "011101101",
                        b"001_0010_000_0110_000_0000" when "011101110",
                        b"001_0010_000_0110_000_0100" when "011101111",

                        b"001_0010_100_1100_000_0001" when "011110000",
                        b"001_0010_100_1100_100_1111" when "011110001",
                        b"001_0010_100_1100_001_0010" when "011110010",
                        b"001_0010_100_1100_000_0110" when "011110011",
                        b"001_0010_100_1100_100_1100" when "011110100",
                        b"001_0010_100_1100_010_0100" when "011110101",
                        b"001_0010_100_1100_010_0000" when "011110110",
                        b"001_0010_100_1100_000_1111" when "011110111",
                        b"001_0010_100_1100_000_0000" when "011111000",
                        b"001_0010_100_1100_000_0100" when "011111001",

                        b"001_0010_010_0100_000_0001" when "011111010",
                        b"001_0010_010_0100_100_1111" when "011111011",
                        b"001_0010_010_0100_001_0010" when "011111100",
                        b"001_0010_010_0100_000_0110" when "011111101",
                        b"001_0010_010_0100_100_1100" when "011111110",
                        b"001_0010_010_0100_010_0100" when "011111111",
                        b"001_0010_010_0100_010_0000" when "100000000",
                        b"001_0010_010_0100_000_1111" when "100000001",
                        b"001_0010_010_0100_000_0000" when "100000010",
                        b"001_0010_010_0100_000_0100" when "100000011",

                        b"001_0010_010_0000_000_0001" when "100000100",
                        b"001_0010_010_0000_100_1111" when "100000101",
                        b"001_0010_010_0000_001_0010" when "100000110",
                        b"001_0010_010_0000_000_0110" when "100000111",
                        b"001_0010_010_0000_100_1100" when "100001000",
                        b"001_0010_010_0000_010_0100" when "100001001",
                        b"001_0010_010_0000_010_0000" when "100001010",
                        b"001_0010_010_0000_000_1111" when "100001011",
                        b"001_0010_010_0000_000_0000" when "100001100",
                        b"001_0010_010_0000_000_0100" when "100001101",

                        b"001_0010_000_1111_000_0001" when "100001110",
                        b"001_0010_000_1111_100_1111" when "100001111",
                        b"001_0010_000_1111_001_0010" when "100010000",
                        b"001_0010_000_1111_000_0110" when "100010001",
                        b"001_0010_000_1111_100_1100" when "100010010",
                        b"001_0010_000_1111_010_0100" when "100010011",
                        b"001_0010_000_1111_010_0000" when "100010100",
                        b"001_0010_000_1111_000_1111" when "100010101",
                        b"001_0010_000_1111_000_0000" when "100010110",
                        b"001_0010_000_1111_000_0100" when "100010111",

                        b"001_0010_000_0000_000_0001" when "100011000",
                        b"001_0010_000_0000_100_1111" when "100011001",
                        b"001_0010_000_0000_001_0010" when "100011010",
                        b"001_0010_000_0000_000_0110" when "100011011",
                        b"001_0010_000_0000_100_1100" when "100011100",
                        b"001_0010_000_0000_010_0100" when "100011101",
                        b"001_0010_000_0000_010_0000" when "100011110",
                        b"001_0010_000_0000_000_1111" when "100011111",
                        b"001_0010_000_0000_000_0000" when "100100000",
                        b"001_0010_000_0000_000_0100" when "100100001",

                        b"001_0010_000_0100_000_0001" when "100100010",
                        b"001_0010_000_0100_100_1111" when "100100011",
                        b"001_0010_000_0100_001_0010" when "100100100",
                        b"001_0010_000_0100_000_0110" when "100100101",
                        b"001_0010_000_0100_100_1100" when "100100110",
                        b"001_0010_000_0100_010_0100" when "100100111",
                        b"001_0010_000_0100_010_0000" when "100101000",
                        b"001_0010_000_0100_000_1111" when "100101001",
                        b"001_0010_000_0100_000_0000" when "100101010",
                        b"001_0010_000_0100_000_0100" when "100101011",

                        b"000_0110_000_0001_000_0001" when "100101100",
                        b"000_0110_000_0001_100_1111" when "100101101",
                        b"000_0110_000_0001_001_0010" when "100101110",
                        b"000_0110_000_0001_000_0110" when "100101111",
                        b"000_0110_000_0001_100_1100" when "100110000",
                        b"000_0110_000_0001_010_0100" when "100110001",
                        b"000_0110_000_0001_010_0000" when "100110010",
                        b"000_0110_000_0001_000_1111" when "100110011",
                        b"000_0110_000_0001_000_0000" when "100110100",
                        b"000_0110_000_0001_000_0100" when "100110101",

                        b"000_0110_100_1111_000_0001" when "100110110",
                        b"000_0110_100_1111_100_1111" when "100110111",
                        b"000_0110_100_1111_001_0010" when "100111000",
                        b"000_0110_100_1111_000_0110" when "100111001",
                        b"000_0110_100_1111_100_1100" when "100111010",
                        b"000_0110_100_1111_010_0100" when "100111011",
                        b"000_0110_100_1111_010_0000" when "100111100",
                        b"000_0110_100_1111_000_1111" when "100111101",
                        b"000_0110_100_1111_000_0000" when "100111110",
                        b"000_0110_100_1111_000_0100" when "100111111",

                        b"000_0110_001_0010_000_0001" when "101000000",
                        b"000_0110_001_0010_100_1111" when "101000001",
                        b"000_0110_001_0010_001_0010" when "101000010",
                        b"000_0110_001_0010_000_0110" when "101000011",
                        b"000_0110_001_0010_100_1100" when "101000100",
                        b"000_0110_001_0010_010_0100" when "101000101",
                        b"000_0110_001_0010_010_0000" when "101000110",
                        b"000_0110_001_0010_000_1111" when "101000111",
                        b"000_0110_001_0010_000_0000" when "101001000",
                        b"000_0110_001_0010_000_0100" when "101001001",

                        b"000_0110_000_0110_000_0001" when "101001010",
                        b"000_0110_000_0110_100_1111" when "101001011",
                        b"000_0110_000_0110_001_0010" when "101001100",
                        b"000_0110_000_0110_000_0110" when "101001101",
                        b"000_0110_000_0110_100_1100" when "101001110",
                        b"000_0110_000_0110_010_0100" when "101001111",
                        b"000_0110_000_0110_010_0000" when "101010000",
                        b"000_0110_000_0110_000_1111" when "101010001",
                        b"000_0110_000_0110_000_0000" when "101010010",
                        b"000_0110_000_0110_000_0100" when "101010011",

                        b"000_0110_100_1100_000_0001" when "101010100",
                        b"000_0110_100_1100_100_1111" when "101010101",
                        b"000_0110_100_1100_001_0010" when "101010110",
                        b"000_0110_100_1100_000_0110" when "101010111",
                        b"000_0110_100_1100_100_1100" when "101011000",
                        b"000_0110_100_1100_010_0100" when "101011001",
                        b"000_0110_100_1100_010_0000" when "101011010",
                        b"000_0110_100_1100_000_1111" when "101011011",
                        b"000_0110_100_1100_000_0000" when "101011100",
                        b"000_0110_100_1100_000_0100" when "101011101",

                        b"000_0110_010_0100_000_0001" when "101011110",
                        b"000_0110_010_0100_100_1111" when "101011111",
                        b"000_0110_010_0100_001_0010" when "101100000",
                        b"000_0110_010_0100_000_0110" when "101100001",
                        b"000_0110_010_0100_100_1100" when "101100010",
                        b"000_0110_010_0100_010_0100" when "101100011",
                        b"000_0110_010_0100_010_0000" when "101100100",
                        b"000_0110_010_0100_000_1111" when "101100101",
                        b"000_0110_010_0100_000_0000" when "101100110",
                        b"000_0110_010_0100_000_0100" when "101100111",

                        b"000_0110_010_0000_000_0001" when "101101000",
                        b"000_0110_010_0000_100_1111" when "101101001",
                        b"000_0110_010_0000_001_0010" when "101101010",
                        b"000_0110_010_0000_000_0110" when "101101011",
                        b"000_0110_010_0000_100_1100" when "101101100",
                        b"000_0110_010_0000_010_0100" when "101101101",
                        b"000_0110_010_0000_010_0000" when "101101110",
                        b"000_0110_010_0000_000_1111" when "101101111",
                        b"000_0110_010_0000_000_0000" when "101110000",
                        b"000_0110_010_0000_000_0100" when "101110001",

                        b"000_0110_000_1111_000_0001" when "101110010",
                        b"000_0110_000_1111_100_1111" when "101110011",
                        b"000_0110_000_1111_001_0010" when "101110100",
                        b"000_0110_000_1111_000_0110" when "101110101",
                        b"000_0110_000_1111_100_1100" when "101110110",
                        b"000_0110_000_1111_010_0100" when "101110111",
                        b"000_0110_000_1111_010_0000" when "101111000",
                        b"000_0110_000_1111_000_1111" when "101111001",
                        b"000_0110_000_1111_000_0000" when "101111010",
                        b"000_0110_000_1111_000_0100" when "101111011",

                        b"000_0110_000_0000_000_0001" when "101111100",
                        b"000_0110_000_0000_100_1111" when "101111101",
                        b"000_0110_000_0000_001_0010" when "101111110",
                        b"000_0110_000_0000_000_0110" when "101111111",
                        b"000_0110_000_0000_100_1100" when "110000000",
                        b"000_0110_000_0000_010_0100" when "110000001",
                        b"000_0110_000_0000_010_0000" when "110000010",
                        b"000_0110_000_0000_000_1111" when "110000011",
                        b"000_0110_000_0000_000_0000" when "110000100",
                        b"000_0110_000_0000_000_0100" when "110000101",

                        b"000_0110_000_0100_000_0001" when "110000110",
                        b"000_0110_000_0100_100_1111" when "110000111",
                        b"000_0110_000_0100_001_0010" when "110001000",
                        b"000_0110_000_0100_000_0110" when "110001001",
                        b"000_0110_000_0100_100_1100" when "110001010",
                        b"000_0110_000_0100_010_0100" when "110001011",
                        b"000_0110_000_0100_010_0000" when "110001100",
                        b"000_0110_000_0100_000_1111" when "110001101",
                        b"000_0110_000_0100_000_0000" when "110001110",
                        b"000_0110_000_0100_000_0100" when "110001111",

                        b"100_1100_000_0001_000_0001" when "110010000",
                        b"100_1100_000_0001_100_1111" when "110010001",
                        b"100_1100_000_0001_001_0010" when "110010010",
                        b"100_1100_000_0001_000_0110" when "110010011",
                        b"100_1100_000_0001_100_1100" when "110010100",
                        b"100_1100_000_0001_010_0100" when "110010101",
                        b"100_1100_000_0001_010_0000" when "110010110",
                        b"100_1100_000_0001_000_1111" when "110010111",
                        b"100_1100_000_0001_000_0000" when "110011000",
                        b"100_1100_000_0001_000_0100" when "110011001",

                        b"100_1100_100_1111_000_0001" when "110011010",
                        b"100_1100_100_1111_100_1111" when "110011011",
                        b"100_1100_100_1111_001_0010" when "110011100",
                        b"100_1100_100_1111_000_0110" when "110011101",
                        b"100_1100_100_1111_100_1100" when "110011110",
                        b"100_1100_100_1111_010_0100" when "110011111",
                        b"100_1100_100_1111_010_0000" when "110100000",
                        b"100_1100_100_1111_000_1111" when "110100001",
                        b"100_1100_100_1111_000_0000" when "110100010",
                        b"100_1100_100_1111_000_0100" when "110100011",

                        b"100_1100_001_0010_000_0001" when "110100100",
                        b"100_1100_001_0010_100_1111" when "110100101",
                        b"100_1100_001_0010_001_0010" when "110100110",
                        b"100_1100_001_0010_000_0110" when "110100111",
                        b"100_1100_001_0010_100_1100" when "110101000",
                        b"100_1100_001_0010_010_0100" when "110101001",
                        b"100_1100_001_0010_010_0000" when "110101010",
                        b"100_1100_001_0010_000_1111" when "110101011",
                        b"100_1100_001_0010_000_0000" when "110101100",
                        b"100_1100_001_0010_000_0100" when "110101101",

                        b"100_1100_000_0110_000_0001" when "110101110",
                        b"100_1100_000_0110_100_1111" when "110101111",
                        b"100_1100_000_0110_001_0010" when "110110000",
                        b"100_1100_000_0110_000_0110" when "110110001",
                        b"100_1100_000_0110_100_1100" when "110110010",
                        b"100_1100_000_0110_010_0100" when "110110011",
                        b"100_1100_000_0110_010_0000" when "110110100",
                        b"100_1100_000_0110_000_1111" when "110110101",
                        b"100_1100_000_0110_000_0000" when "110110110",
                        b"100_1100_000_0110_000_0100" when "110110111",

                        b"100_1100_100_1100_000_0001" when "110111000",
                        b"100_1100_100_1100_100_1111" when "110111001",
                        b"100_1100_100_1100_001_0010" when "110111010",
                        b"100_1100_100_1100_000_0110" when "110111011",
                        b"100_1100_100_1100_100_1100" when "110111100",
                        b"100_1100_100_1100_010_0100" when "110111101",
                        b"100_1100_100_1100_010_0000" when "110111110",
                        b"100_1100_100_1100_000_1111" when "110111111",
                        b"100_1100_100_1100_000_0000" when "111000000",
                        b"100_1100_100_1100_000_0100" when "111000001",

                        b"100_1100_010_0100_000_0001" when "111000010",
                        b"100_1100_010_0100_100_1111" when "111000011",
                        b"100_1100_010_0100_001_0010" when "111000100",
                        b"100_1100_010_0100_000_0110" when "111000101",
                        b"100_1100_010_0100_100_1100" when "111000110",
                        b"100_1100_010_0100_010_0100" when "111000111",
                        b"100_1100_010_0100_010_0000" when "111001000",
                        b"100_1100_010_0100_000_1111" when "111001001",
                        b"100_1100_010_0100_000_0000" when "111001010",
                        b"100_1100_010_0100_000_0100" when "111001011",

                        b"100_1100_010_0000_000_0001" when "111001100",
                        b"100_1100_010_0000_100_1111" when "111001101",
                        b"100_1100_010_0000_001_0010" when "111001110",
                        b"100_1100_010_0000_000_0110" when "111001111",
                        b"100_1100_010_0000_100_1100" when "111010000",
                        b"100_1100_010_0000_010_0100" when "111010001",
                        b"100_1100_010_0000_010_0000" when "111010010",
                        b"100_1100_010_0000_000_1111" when "111010011",
                        b"100_1100_010_0000_000_0000" when "111010100",
                        b"100_1100_010_0000_000_0100" when "111010101",

                        b"100_1100_000_1111_000_0001" when "111010110",
                        b"100_1100_000_1111_100_1111" when "111010111",
                        b"100_1100_000_1111_001_0010" when "111011000",
                        b"100_1100_000_1111_000_0110" when "111011001",
                        b"100_1100_000_1111_100_1100" when "111011010",
                        b"100_1100_000_1111_010_0100" when "111011011",
                        b"100_1100_000_1111_010_0000" when "111011100",
                        b"100_1100_000_1111_000_1111" when "111011101",
                        b"100_1100_000_1111_000_0000" when "111011110",
                        b"100_1100_000_1111_000_0100" when "111011111",

                        b"100_1100_000_0000_000_0001" when "111100000",
                        b"100_1100_000_0000_100_1111" when "111100001",
                        b"100_1100_000_0000_001_0010" when "111100010",
                        b"100_1100_000_0000_000_0110" when "111100011",
                        b"100_1100_000_0000_100_1100" when "111100100",
                        b"100_1100_000_0000_010_0100" when "111100101",
                        b"100_1100_000_0000_010_0000" when "111100110",
                        b"100_1100_000_0000_000_1111" when "111100111",
                        b"100_1100_000_0000_000_0000" when "111101000",
                        b"100_1100_000_0000_000_0100" when "111101001",

                        b"100_1100_000_0100_000_0001" when "111101010",
                        b"100_1100_000_0100_100_1111" when "111101011",
                        b"100_1100_000_0100_001_0010" when "111101100",
                        b"100_1100_000_0100_000_0110" when "111101101",
                        b"100_1100_000_0100_100_1100" when "111101110",
                        b"100_1100_000_0100_010_0100" when "111101111",
                        b"100_1100_000_0100_010_0000" when "111110000",
                        b"100_1100_000_0100_000_1111" when "111110001",
                        b"100_1100_000_0100_000_0000" when "111110010",
                        b"100_1100_000_0100_000_0100" when "111110011",

                        b"010_0100_000_0001_000_0001" when "111110100",
                        b"010_0100_000_0001_100_1111" when "111110101",
                        b"010_0100_000_0001_001_0010" when "111110110",
                        b"010_0100_000_0001_000_0110" when "111110111",

                        b"000_0000_000_0000_000_0000" when others;

                        
end Behavioral;